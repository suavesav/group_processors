`include "pipeline_register_if.vh"

module ifid
  import cpu_types_pkg::*;
  (
    input logic CLK, nRST,
    pipeline_register_if.ifid ifidif
  );

  always_ff @(posedge CLK, negedge nRST)
  begin
    if (!nRST)
    begin
    end
    else if(ifidif.ifW)
    begin
    end
  end
endmodule // FETCH_DECODE
