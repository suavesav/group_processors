`include "hazard_unit_if.vh"
`include "cpu_types_pkg.vh"
