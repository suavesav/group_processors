//`include "cache_control_if.vh"
//`include "datapath_cache_if.vh"

module ICACHE(
	      input cache_control_if.cc ccif,
	      input datapath_cache_if.dc dcif
	      );

   
